package uart_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import wb_agt_pkg::*;
  `include "uart_env_config.sv"
  `include "uart_scoreboard.sv"
  `include "uart_env.sv"
endpackage